library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity MemoryManager is
	port (
		clk : in std_logic;
		efm_mode : in boolean;
		ebi_data : in std_logic_vector(15 downto 0)
end MemoryManager;

architecture Behavioral of MemoryManager is

begin


end Behavioral;

